module alu(
  // 演算対象
  input [15:0] a,
  input [15:0] b,

  // 操作コード
  input [3:0] op,

  // 演算結果
  output reg [15:0] res,

  // 条件コード
  output reg [3:0] szcv);

  // 右算術シフトのために符号ありのb[3:0]を保持するレジスタ
  reg signed [3:0] bb;

  // 桁上げを保持するレジスタ
  reg carry;


  // シフトを行う関数
  function [16:0] shift;
  input [3:0] opcode;
  begin
    if(opcode == 4'b1000) begin
      // 左論理シフト（空いた部分は0で埋める）
      case (b[3:0])
      4'b0000: shift = {1'b0,a[15:0]};
      4'b0001: shift = {a[15:0],1'b0};
      4'b0010: shift = {a[14:0],2'b00};
      4'b0011: shift = {a[13:0],3'b000};
      4'b0100: shift = {a[12:0],4'b0000};
      4'b0101: shift = {a[11:0],5'b00000};
      4'b0110: shift = {a[10:0],6'b000000};
      4'b0111: shift = {a[9:0],7'b0000000};
      4'b1000: shift = {a[8:0],8'b00000000};
      4'b1001: shift = {a[7:0],9'b000000000};
      4'b1010: shift = {a[6:0],10'b0000000000};
      4'b1011: shift = {a[5:0],11'b00000000000};
      4'b1100: shift = {a[4:0],12'b000000000000};
      4'b1101: shift = {a[3:0],13'b0000000000000};
      4'b1110: shift = {a[2:0],14'b00000000000000};
      4'b1111: shift = {a[1:0],15'b000000000000000};
      default: shift = 16'b0000_0000_0000_0000;
      endcase
    end
    else if(opcode == 4'b1001) begin
      // 左循環シフト（空いた部分はシフトアウトされたビット列）
      case (b[3:0])
      4'b0000: shift = {1'b0,a[15:0]};
      4'b0001: shift = {1'b0,a[14:0],a[15]};
      4'b0010: shift = {1'b0,a[13:0],a[15:14]};
      4'b0011: shift = {1'b0,a[12:0],a[15:13]};
      4'b0100: shift = {1'b0,a[11:0],a[15:12]};
      4'b0101: shift = {1'b0,a[10:0],a[15:11]};
      4'b0110: shift = {1'b0,a[9:0],a[15:10]};
      4'b0111: shift = {1'b0,a[8:0],a[15:9]};
      4'b1000: shift = {1'b0,a[7:0],a[15:8]};
      4'b1001: shift = {1'b0,a[6:0],a[15:7]};
      4'b1010: shift = {1'b0,a[5:0],a[15:6]};
      4'b1011: shift = {1'b0,a[4:0],a[15:5]};
      4'b1100: shift = {1'b0,a[3:0],a[15:4]};
      4'b1101: shift = {1'b0,a[2:0],a[15:3]};
      4'b1110: shift = {1'b0,a[1:0],a[15:2]};
      4'b1111: shift = {1'b0,a[0],a[15:1]};
      default: shift = {1'b0,16'b0000_0000_0000_0000};
      endcase
    end
    else if(opcode == 4'b1010) begin
      // 右論理シフト（空いた部分は0で埋める）
      case (b[3:0])
      4'b0000: shift = {1'b0,a[15:0]};
      4'b0001: shift = {a[0],1'b0,a[15:1]};
      4'b0010: shift = {a[1],2'b00,a[15:2]};
      4'b0011: shift = {a[2],3'b000,a[15:3]};
      4'b0100: shift = {a[3],4'b0000,a[15:4]};
      4'b0101: shift = {a[4],5'b00000,a[15:5]};
      4'b0110: shift = {a[5],6'b000000,a[15:6]};
      4'b0111: shift = {a[6],7'b0000000,a[15:7]};
      4'b1000: shift = {a[7],8'b00000000,a[15:8]};
      4'b1001: shift = {a[8],9'b000000000,a[15:9]};
      4'b1010: shift = {a[9],10'b0000000000,a[15:10]};
      4'b1011: shift = {a[10],11'b00000000000,a[15:11]};
      4'b1100: shift = {a[11],12'b000000000000,a[15:12]};
      4'b1101: shift = {a[12],13'b0000000000000,a[15:13]};
      4'b1110: shift = {a[13],14'b00000000000000,a[15:14]};
      4'b1111: shift = {a[14],15'b000000000000000,a[15]};
      default: shift = {1'b0,16'b0000_0000_0000_0000};
      endcase
    end
    else if(opcode == 4'b1011) begin
      // 右算術シフト（空いた部分は符号ビットで埋める）
      if(a[15] == 1'b0) begin
        //符号ビットが0
        case (b[3:0])
        4'b0000: shift = {1'b0,a[15:0]};
        4'b0001: shift = {a[0],1'b0,a[15:1]};
        4'b0010: shift = {a[1],2'b00,a[15:2]};
        4'b0011: shift = {a[2],3'b000,a[15:3]};
        4'b0100: shift = {a[3],4'b0000,a[15:4]};
        4'b0101: shift = {a[4],5'b00000,a[15:5]};
        4'b0110: shift = {a[5],6'b000000,a[15:6]};
        4'b0111: shift = {a[6],7'b0000000,a[15:7]};
        4'b1000: shift = {a[7],8'b00000000,a[15:8]};
        4'b1001: shift = {a[8],9'b000000000,a[15:9]};
        4'b1010: shift = {a[9],10'b0000000000,a[15:10]};
        4'b1011: shift = {a[10],11'b00000000000,a[15:11]};
        4'b1100: shift = {a[11],12'b000000000000,a[15:12]};
        4'b1101: shift = {a[12],13'b0000000000000,a[15:13]};
        4'b1110: shift = {a[13],14'b00000000000000,a[15:14]};
        4'b1111: shift = {a[14],15'b000000000000000,a[15]};
        default: shift = {1'b0,16'b0000_0000_0000_0000};
        endcase
      end
      else begin
        // 符号ビットが1
        case(b[3:0])
        4'b0000: shift = {1'b0,a[15:0]};
        4'b0001: shift = {a[0],1'b1,a[15:1]};
        4'b0010: shift = {a[1],2'b11,a[15:3]};
        4'b0100: shift = {a[3],4'b1111,a[15:4]};
        4'b0101: shift = {a[4],5'b11111,a[15:5]};
        4'b0110: shift = {a[5],6'b111111,a[15:6]};
        4'b0111: shift = {a[6],7'b1111111,a[15:7]};
        4'b1000: shift = {a[7],8'b11111111,a[15:8]};
        4'b1001: shift = {a[8],9'b111111111,a[15:9]};
        4'b1010: shift = {a[9],10'b1111111111,a[15:10]};
        4'b1011: shift = {a[10],11'b11111111111,a[15:11]};
        4'b1100: shift = {a[11],12'b111111111111,a[15:12]};
        4'b1101: shift = {a[12],13'b1111111111111,a[15:13]};
        4'b1110: shift = {a[13],14'b11111111111111,a[15:14]};
        4'b1111: shift = {a[14],15'b111111111111111,a[15]};
        default: shift = {1'b0,16'b0000_0000_0000_0000};
        endcase
      end
    end 
    else begin
      //操作コードがシフト演算ではないとき
      shift = {1'b0,16'b0000_0000_0000_0000};
    end
  end
  endfunction

  always @* begin
    bb <= b[3:0];
    case(op)
    4'b0000: {carry,res} <= a + b;
    4'b0001: {carry,res} <= a - b;
    4'b0010: {carry,res} <= {1'b0,a & b};
    4'b0011: {carry,res} <= {1'b0,a | b};
    4'b0100: {carry,res} <= {1'b0,a ^ b};
    4'b0101: {carry,res} <= a - b;
    4'b0110: {carry,res} <= {1'b0,b[15:0]};
    4'b1000: {carry,res} <= shift(op);
    4'b1001: {carry,res} <= shift(op);        
    4'b1010: {carry,res} <= shift(op);
    4'b1011: {carry,res} <= shift(op);
    default: {carry,res} <= {1'b0,16'b0000_0000_0000_0000};	 
    endcase

    // 正負のフラグ
    szcv[3] <= res[15];

    // ゼロかどうかのフラグ
    if(res == 16'b0000_0000_0000_0000) begin
      szcv[2] = 1'b1;
    end
    else begin
      szcv[2] = 1'b0;
    end
    
    // 桁上げのフラグ
    szcv[1] <= carry;

    // オーバーフローのフラグ
    if(op == 4'b0000 && a[15] == b[15] && a[15] != res[15]) begin
      szcv[0] = 1'b1;
    end
    else if(op == 4'b0001 && a[15] == res[15] && a[15] != b[15]) begin
      szcv[0] = 1'b1;
    end
    else begin
      szcv[0] = 1'b0;
    end

  end

endmodule