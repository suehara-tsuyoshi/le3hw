module chattering(
  input clock,
  input reset,
  input exec,
  output reg state);

  reg [31:0] time_counter = 32'b0000_0000_0000_0000_0000_0000_0000_0000;

  always @(posedge clock) begin
    if(reset == 1'b0) begin
      time_counter <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
      state <= 1'b0;
    end
    else if(exec == 1'b0) begin
      time_counter <= time_counter + 1;
      if(time_counter == 32'b0000_0000_0000_0010_0000_0000_0000_0000) begin
        if(state == 1'b0) begin
          state <= 1'b1;
        end 
        else if(state == 1'b1) begin
          state <= 1'b0;
        end
      end
    end
    else begin
      time_counter <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
      state <= state;
    end
  end
endmodule